-------------------------------------------------------------------------------
--
-- Title       : TutorVHDL
-- Design      : TutorVHDL
-- Author      : J.Kasperek & P.J.Rajda
-- Company     : AGH Krak�w
--
-------------------------------------------------------------------------------
--
-- Description : 
-- Synchronous 3bits binary up counter with synchronous reset
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity TutorVHDL is
port (
   clk: in std_logic; -- 100MHz clock input 
   DUTY_INCREASE: in std_logic; -- button to increase duty cycle by 10%
   DUTY_DECREASE: in std_logic; -- button to decrease duty cycle by 10%
   PWM_OUT: out std_logic -- PWM signal out with frequency of 10MHz
  );
end TutorVHDL;

architecture Behavioral of TutorVHDL is
 -- D-Flip-Flop for debouncing module
 component Debouncer   --DFF Debunce
 Port ( 
  CLK : in std_logic;
  en : in std_logic;
  D : in std_logic;
  Q : out std_logic
  );
 end component;
 signal slow_clk_en: std_logic:='0'; -- slow clock enable for debouncing
 signal counter_slow: std_logic_vector(27 downto 0):=(others => '0');-- counter for creating slow clock
 signal tmp1,tmp2,duty_inc: std_logic;-- temporary signals for deboucing
 signal tmp3,tmp4,duty_dec: std_logic;-- temporary signals for deboucing
 signal counter_PWM: std_logic_vector(3 downto 0):=(others => '0');-- counter for PWM signal
 signal DUTY_CYCLE: std_logic_vector(3 downto 0):=x"5";
begin
 -- Debouncing process
 -- First generate slow clock enable for deboucing (4Hz)
 process(clk)
 begin
  if(rising_edge(clk)) then
   counter_slow <= counter_slow + x"0000001";
   --if(counter_slow>=x"17D7840") then -- for running on FPGA -- comment when running simulation
   if(counter_slow>=x"0000001") then -- for running simulation -- comment when running on FPGA
    counter_slow <= x"0000000";
   end if;
  end if;
 end process;
 --slow_clk_en <= '1' when counter_slow = x"17D7840" else '0';-- for running on FPGA -- comment when running simulation 
 slow_clk_en <= '1' when counter_slow = x"000001" else '0';-- for running simulation -- comment when running on FPGA
 -- debounce part for duty increasing button
 stage0: Debouncer port map(clk,slow_clk_en , DUTY_INCREASE, tmp1);
 stage1: Debouncer port map(clk,slow_clk_en , tmp1, tmp2); 
 duty_inc <=  tmp1 and (not tmp2) and slow_clk_en;
 -- debounce part for duty decreasing button
 stage2: Debouncer port map(clk,slow_clk_en , DUTY_DECREASE, tmp3);
 stage3: Debouncer port map(clk,slow_clk_en , tmp3, tmp4); 
 duty_dec <=  tmp3 and (not tmp4) and slow_clk_en;
 -- for controlling duty cycle by these buttons
 process(clk)
 begin
  if(rising_edge(clk)) then
   if(duty_inc='1' and DUTY_CYCLE <= x"9") then
    DUTY_CYCLE <= DUTY_CYCLE + x"1";--increase duty cycle by 10%
   elsif(duty_dec='1' and DUTY_CYCLE>=x"1") then
    DUTY_CYCLE <= DUTY_CYCLE - x"1";--decrease duty cycle by 10%
   end if;
  end if;
 end process;
 -- Create 10MHz PWM signal
 process(clk)
 begin
  if(rising_edge(clk)) then
   counter_PWM <= counter_PWM + x"1";
   if(counter_PWM>=x"9") then
    counter_PWM <= x"0";
   end if;
  end if;
 end process;
 PWM_OUT <= '1' when counter_PWM < DUTY_CYCLE else '0';
end Behavioral;