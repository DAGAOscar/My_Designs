//-----------------------------------------------------------------------------
//
// Title       : tutorvhdl_tb_tim
// Design      : TutorVHDL
// Author      : IE
// Company     : AGH
//
//-----------------------------------------------------------------------------
//
// File        : TutorVHDL_TB.v
// Generated   : Wed Dec  8 10:45:16 2021
// From        : C:\My_Designs\Tutorials_cz0940_LF\TutorVHDL_Sr0940\src\tutorvhdl_TB_tim\TutorVHDL_TB_settings.txt
// By          : tb_verilog.pl ver. ver 1.2s
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------

`timescale 1ps / 1ps
module tutorvhdl_tb_tim;


//Internal signals declarations:
reg CLR;
reg CLK;
reg CE;
reg LOAD;
reg DIR;
reg SEL;
reg [3:0]DATA;
reg OE;
reg LE;
wire [3:0]Q;



// Unit Under Test port map
	TutorVHDL UUT (
		.CLR(CLR),
		.CLK(CLK),
		.CE(CE),
		.LOAD(LOAD),
		.DIR(DIR),
		.SEL(SEL),
		.DATA(DATA),
		.OE(OE),
		.LE(LE),
		.Q(Q));

initial
	$monitor($realtime,,"ps %h %h %h %h %h %h %h %h %h %h ",CLR,CLK,CE,LOAD,DIR,SEL,DATA,OE,LE,Q);

//Below code was generated based on waveform file: "C:\My_Designs\Tutorials_cz0940_LF\TutorVHDL_Sr0940\compile\TutorVHDL.ver"

initial
begin : STIMUL // begin of stimulus process
	#0
	CE = 1'b1;
	LOAD = 1'b0;
	SEL = 1'b0;
	CLR = 1'b0;
	DIR = 1'b1;
	CLK = 1'b0;
	LE = 1'b0;
	OE = 1'b1;
	DATA = 4'b0110;
    #50000; //0
	CLK = 1'b1;
    #25000; //50000
	CLR = 1'b1;
    #25000; //75000
	CLK = 1'b0;
    #50000; //100000
	CLK = 1'b1;
    #25000; //150000
	CLR = 1'b0;
    #25000; //175000
	CLK = 1'b0;
    #50000; //200000
	CLK = 1'b1;
    #50000; //250000
	LOAD = 1'b1;
	CLK = 1'b0;
    #50000; //300000
	CLK = 1'b1;
    #50000; //350000
	CLK = 1'b0;
    #50000; //400000
	CLK = 1'b1;
    #50000; //450000
	LOAD = 1'b0;
	CLK = 1'b0;
    #50000; //500000
	CLK = 1'b1;
    #50000; //550000
	CLK = 1'b0;
    #50000; //600000
	CLK = 1'b1;
    #50000; //650000
	CLK = 1'b0;
    #50000; //700000
	CLK = 1'b1;
    #50000; //750000
	CLK = 1'b0;
    #50000; //800000
	CLK = 1'b1;
    #50000; //850000
	CLK = 1'b0;
    #50000; //900000
	CLK = 1'b1;
    #50000; //950000
	CE = 1'b0;
	CLK = 1'b0;
    #50000; //1000000
	CLK = 1'b1;
    #50000; //1050000
	CLK = 1'b0;
    #50000; //1100000
	CLK = 1'b1;
    #50000; //1150000
	CLK = 1'b0;
    #50000; //1200000
	CLK = 1'b1;
    #50000; //1250000
	CE = 1'b1;
	CLK = 1'b0;
    #50000; //1300000
	CLK = 1'b1;
    #50000; //1350000
	DIR = 1'b0;
	CLK = 1'b0;
    #50000; //1400000
	CLK = 1'b1;
    #50000; //1450000
	CLK = 1'b0;
    #50000; //1500000
	CLK = 1'b1;
    #50000; //1550000
	CLK = 1'b0;
    #50000; //1600000
	CLK = 1'b1;
    #50000; //1650000
	CLK = 1'b0;
    #50000; //1700000
	CLK = 1'b1;
    #50000; //1750000
	CLK = 1'b0;
    #50000; //1800000
	CLK = 1'b1;
    #50000; //1850000
	CLK = 1'b0;
    #50000; //1900000
	CLK = 1'b1;
    #50000; //1950000
	CLK = 1'b0;
    #50000; //2000000
	CLK = 1'b1;
    #50000; //2050000
	CLK = 1'b0;
    #50000; //2100000
	CLK = 1'b1;
    #50000; //2150000
	CLK = 1'b0;
    #50000; //2200000
	CLK = 1'b1;
    #50000; //2250000
	CLK = 1'b0;
    #50000; //2300000
	CLK = 1'b1;
    #50000; //2350000
	CLK = 1'b0;
    #50000; //2400000
	CLK = 1'b1;
    #50000; //2450000
	CLK = 1'b0;
	OE = 1'b0;
    #50000; //2500000
	CLK = 1'b1;
    #50000; //2550000
	CLK = 1'b0;
	OE = 1'b1;
    #50000; //2600000
	CLK = 1'b1;
    #25000; //2650000
	CLR = 1'b1;
    #25000; //2675000
	CLK = 1'b0;
    #50000; //2700000
	CLK = 1'b1;
    #50000; //2750000
	CLK = 1'b0;
    #50000; //2800000
	CLK = 1'b1;
    #25000; //2850000
	CLR = 1'b0;
    #25000; //2875000
	CLK = 1'b0;
    #50000; //2900000
	CLK = 1'b1;
    #50000; //2950000
	SEL = 1'b1;
	CLK = 1'b0;
    #50000; //3000000
	CLK = 1'b1;
    #50000; //3050000
	CLK = 1'b0;
    #50000; //3100000
	CLK = 1'b1;
    #50000; //3150000
	CLK = 1'b0;
    #50000; //3200000
	CLK = 1'b1;
	LE = 1'b1;
    #50000; //3250000
	CLK = 1'b0;
    #50000; //3300000
	CLK = 1'b1;
	DATA = 4'b0001;
    #50000; //3350000
	CLK = 1'b0;
    #50000; //3400000
	CLK = 1'b1;
	LE = 1'b0;
    #50000; //3450000
	CLK = 1'b0;
    #50000; //3500000
	CLK = 1'b1;
	DATA = 4'b0101;
    #50000; //3550000
	CLK = 1'b0;
    #50000; //3600000
	CLK = 1'b1;
    #50000; //3650000
	CLK = 1'b0;
    #50000; //3700000
	CLK = 1'b1;
    #50000; //3750000
	SEL = 1'b0;
	CLK = 1'b0;
    #50000; //3800000
	CLK = 1'b1;
    #50000; //3850000
	CLK = 1'b0;
    #50000; //3900000
	CLK = 1'b1;
    #50000; //3950000
	CLK = 1'b0;
    #50000; //4000000
	CLK = 1'b1;
    #50000; //4050000
	CLK = 1'b0;
    #50000; //4100000
	CLK = 1'b1;
    #50000; //4150000
	CLK = 1'b0;
    #50000; //4200000
	CLK = 1'b1;
    #50000; //4250000
	CLK = 1'b0;
    #50000; //4300000
	CLK = 1'b1;
    #50000; //4350000
	CLK = 1'b0;
    #50000; //4400000
	CLK = 1'b1;
    #50000; //4450000
	CLK = 1'b0;
    #50000; //4500000
	CLK = 1'b1;
    #50000; //4550000
	CLK = 1'b0;
    #50000; //4600000
	CLK = 1'b1;
    #50000; //4650000
	CLK = 1'b0;
    #50000; //4700000
	CLK = 1'b1;
    #50000; //4750000
	CLK = 1'b0;
    #50000; //4800000
	CLK = 1'b1;
    #50000; //4850000
	CLK = 1'b0;
    #50000; //4900000
	CLK = 1'b1;
    #50000; //4950000
	CLK = 1'b0;
    #50000; //5000000
	CLK = 1'b1;
    #50000; //5050000
	CLK = 1'b0;
    #50000; //5100000
	CLK = 1'b1;
    #50000; //5150000
	CLK = 1'b0;
    #50000; //5200000
	CLK = 1'b1;
    #50000; //5250000
	CLK = 1'b0;
    #50000; //5300000
	CLK = 1'b1;
    #50000; //5350000
	CLK = 1'b0;
    #50000; //5400000
	CLK = 1'b1;
    #50000; //5450000
	CLK = 1'b0;
    #50000; //5500000
	CLK = 1'b1;
    #50000; //5550000
	CLK = 1'b0;
    #50000; //5600000
	CLK = 1'b1;
    #50000; //5650000
	CLK = 1'b0;
    #50000; //5700000
	CLK = 1'b1;
    #50000; //5750000
	CLK = 1'b0;
    #50000; //5800000
	CLK = 1'b1;
    #50000; //5850000
	CLK = 1'b0;
    #50000; //5900000
	CLK = 1'b1;
    #50000; //5950000
	CLK = 1'b0;
end // end of stimulus process
	



endmodule
