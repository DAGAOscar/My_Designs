-------------------------------------------------------------------------------
--
-- Title       : Fub1
-- Design      : TutorVHDL
-- Author      : loueke@student.agh.edu.pl
-- Company     : AGH University of Technology
--
-------------------------------------------------------------------------------
--
-- File        : C:/Users/ferna/Downloads/Tuto_prescaler_LF/TutorVHDL/src/Fub1.vhd
-- Generated   : Tue Dec 21 11:05:39 2021
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Fub1} architecture {Fub1}}



entity Fub1 is
end Fub1;

--}} End of automatically maintained section

architecture Fub1 of Fub1 is
begin

	 -- enter your statements here --

end Fub1;
